
module cx_system (
	altpll_0_locked_conduit_export,
	bme280_i2c_0_control_conduit_busy_out,
	bme280_i2c_0_control_conduit_continuous,
	bme280_i2c_0_control_conduit_enable,
	bme280_i2c_0_i2c_interface_i2c_ack_error,
	bme280_i2c_0_i2c_interface_i2c_addr,
	bme280_i2c_0_i2c_interface_i2c_busy,
	bme280_i2c_0_i2c_interface_i2c_data_rd,
	bme280_i2c_0_i2c_interface_i2c_data_wr,
	bme280_i2c_0_i2c_interface_i2c_ena,
	bme280_i2c_0_i2c_interface_i2c_rw,
	cfg_input_data,
	cfg_input_error,
	cfg_input_valid,
	cfg_output_data,
	cfg_output_error,
	cfg_output_valid,
	clk_clk,
	control_conduit_busy_out,
	fe_ics52000_0_cfg_input_data,
	fe_ics52000_0_cfg_input_error,
	fe_ics52000_0_cfg_input_valid,
	fpga_control_conduit_busy_out,
	fpga_rj45_interface_serial_data_in,
	fpga_rj45_interface_serial_data_out,
	fpga_rj45_interface_serial_clk_out,
	fpga_serial_clk_clk,
	i2c_clk_clk,
	ics52000_physical_mic_data_in,
	ics52000_physical_mic_ws_out,
	ics52000_physical_clk,
	ics52000_physical_mics_rdy,
	led_output_led_sd,
	led_output_led_ws,
	mic_output_channel,
	mic_output_data,
	mic_output_error,
	mic_output_valid,
	ncp5623b_i2c_conduit_i2c_enable_out,
	ncp5623b_i2c_conduit_i2c_address_out,
	ncp5623b_i2c_conduit_i2c_rdwr_out,
	ncp5623b_i2c_conduit_i2c_data_write_out,
	ncp5623b_i2c_conduit_i2c_bsy_in,
	ncp5623b_i2c_conduit_i2c_data_read_in,
	ncp5623b_i2c_conduit_i2c_req_out,
	ncp5623b_i2c_conduit_i2c_rdy_in,
	pll_mclk_clk,
	reset_reset_n,
	rgb_input_data,
	rgb_input_error,
	rgb_input_valid,
	rj45_interface_serial_data_in,
	rj45_interface_serial_data_out,
	serial_clk_clk,
	bme_output_data,
	bme_output_error,
	bme_output_valid);	

	output		altpll_0_locked_conduit_export;
	output		bme280_i2c_0_control_conduit_busy_out;
	input		bme280_i2c_0_control_conduit_continuous;
	input		bme280_i2c_0_control_conduit_enable;
	input		bme280_i2c_0_i2c_interface_i2c_ack_error;
	output	[6:0]	bme280_i2c_0_i2c_interface_i2c_addr;
	input		bme280_i2c_0_i2c_interface_i2c_busy;
	input	[7:0]	bme280_i2c_0_i2c_interface_i2c_data_rd;
	output	[7:0]	bme280_i2c_0_i2c_interface_i2c_data_wr;
	output		bme280_i2c_0_i2c_interface_i2c_ena;
	output		bme280_i2c_0_i2c_interface_i2c_rw;
	input	[15:0]	cfg_input_data;
	input	[1:0]	cfg_input_error;
	input		cfg_input_valid;
	output	[15:0]	cfg_output_data;
	output	[1:0]	cfg_output_error;
	output		cfg_output_valid;
	input		clk_clk;
	output		control_conduit_busy_out;
	input	[15:0]	fe_ics52000_0_cfg_input_data;
	input	[1:0]	fe_ics52000_0_cfg_input_error;
	input		fe_ics52000_0_cfg_input_valid;
	output		fpga_control_conduit_busy_out;
	input		fpga_rj45_interface_serial_data_in;
	output		fpga_rj45_interface_serial_data_out;
	output		fpga_rj45_interface_serial_clk_out;
	input		fpga_serial_clk_clk;
	output		i2c_clk_clk;
	input	[15:0]	ics52000_physical_mic_data_in;
	output	[15:0]	ics52000_physical_mic_ws_out;
	output	[3:0]	ics52000_physical_clk;
	output		ics52000_physical_mics_rdy;
	output		led_output_led_sd;
	output		led_output_led_ws;
	output	[3:0]	mic_output_channel;
	output	[31:0]	mic_output_data;
	output	[1:0]	mic_output_error;
	output		mic_output_valid;
	output		ncp5623b_i2c_conduit_i2c_enable_out;
	output	[6:0]	ncp5623b_i2c_conduit_i2c_address_out;
	output		ncp5623b_i2c_conduit_i2c_rdwr_out;
	output	[7:0]	ncp5623b_i2c_conduit_i2c_data_write_out;
	input		ncp5623b_i2c_conduit_i2c_bsy_in;
	input	[7:0]	ncp5623b_i2c_conduit_i2c_data_read_in;
	output		ncp5623b_i2c_conduit_i2c_req_out;
	input		ncp5623b_i2c_conduit_i2c_rdy_in;
	output		pll_mclk_clk;
	input		reset_reset_n;
	input	[15:0]	rgb_input_data;
	input	[1:0]	rgb_input_error;
	input		rgb_input_valid;
	input		rj45_interface_serial_data_in;
	output		rj45_interface_serial_data_out;
	input		serial_clk_clk;
	output	[95:0]	bme_output_data;
	output	[1:0]	bme_output_error;
	output		bme_output_valid;
endmodule
