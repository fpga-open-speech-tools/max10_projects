-- cx_system.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity cx_system is
	port (
		altpll_0_locked_conduit_export           : out std_logic;                                        --      altpll_0_locked_conduit.export
		bme280_i2c_0_bme_output_data             : out std_logic_vector(95 downto 0);                    --      bme280_i2c_0_bme_output.data
		bme280_i2c_0_bme_output_error            : out std_logic_vector(1 downto 0);                     --                             .error
		bme280_i2c_0_bme_output_valid            : out std_logic;                                        --                             .valid
		bme280_i2c_0_control_conduit_busy_out    : out std_logic;                                        -- bme280_i2c_0_control_conduit.busy_out
		bme280_i2c_0_control_conduit_continuous  : in  std_logic                     := '0';             --                             .continuous
		bme280_i2c_0_control_conduit_enable      : in  std_logic                     := '0';             --                             .enable
		bme280_i2c_0_i2c_interface_i2c_ack_error : in  std_logic                     := '0';             --   bme280_i2c_0_i2c_interface.i2c_ack_error
		bme280_i2c_0_i2c_interface_i2c_addr      : out std_logic_vector(6 downto 0);                     --                             .i2c_addr
		bme280_i2c_0_i2c_interface_i2c_busy      : in  std_logic                     := '0';             --                             .i2c_busy
		bme280_i2c_0_i2c_interface_i2c_data_rd   : in  std_logic_vector(7 downto 0)  := (others => '0'); --                             .i2c_data_rd
		bme280_i2c_0_i2c_interface_i2c_data_wr   : out std_logic_vector(7 downto 0);                     --                             .i2c_data_wr
		bme280_i2c_0_i2c_interface_i2c_ena       : out std_logic;                                        --                             .i2c_ena
		bme280_i2c_0_i2c_interface_i2c_rw        : out std_logic;                                        --                             .i2c_rw
		clk_clk                                  : in  std_logic                     := '0';             --                          clk.clk
		reset_reset_n                            : in  std_logic                     := '0'              --                        reset.reset_n
	);
end entity cx_system;

architecture rtl of cx_system is
	component cx_system_altpll_0 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			locked             : out std_logic;                                        -- export
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			c3                 : out std_logic;                                        -- clk
			c4                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component cx_system_altpll_0;

	component FE_CPLD_BME280_I2C_Reader is
		generic (
			sdo              : std_logic := '0';
			reads_per_second : integer   := 16;
			input_clk        : integer   := 50000000
		);
		port (
			reset_n          : in  std_logic                     := 'X';             -- reset_n
			sys_clk          : in  std_logic                     := 'X';             -- clk
			bme_output_data  : out std_logic_vector(95 downto 0);                    -- data
			bme_output_error : out std_logic_vector(1 downto 0);                     -- error
			bme_output_valid : out std_logic;                                        -- valid
			busy_out         : out std_logic;                                        -- busy_out
			continuous       : in  std_logic                     := 'X';             -- continuous
			enable           : in  std_logic                     := 'X';             -- enable
			i2c_ack_error    : in  std_logic                     := 'X';             -- i2c_ack_error
			i2c_addr         : out std_logic_vector(6 downto 0);                     -- i2c_addr
			i2c_busy         : in  std_logic                     := 'X';             -- i2c_busy
			i2c_data_rd      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- i2c_data_rd
			i2c_data_wr      : out std_logic_vector(7 downto 0);                     -- i2c_data_wr
			i2c_ena          : out std_logic;                                        -- i2c_ena
			i2c_rw           : out std_logic                                         -- i2c_rw
		);
	end component FE_CPLD_BME280_I2C_Reader;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal rst_controller_reset_out_reset           : std_logic; -- rst_controller:reset_out -> [altpll_0:reset, rst_controller_reset_out_reset:in]
	signal reset_reset_n_ports_inv                  : std_logic; -- reset_reset_n:inv -> rst_controller:reset_in0
	signal rst_controller_reset_out_reset_ports_inv : std_logic; -- rst_controller_reset_out_reset:inv -> bme280_i2c_0:reset_n

begin

	altpll_0 : component cx_system_altpll_0
		port map (
			clk                => clk_clk,                        --       inclk_interface.clk
			reset              => rst_controller_reset_out_reset, -- inclk_interface_reset.reset
			read               => open,                           --             pll_slave.read
			write              => open,                           --                      .write
			address            => open,                           --                      .address
			readdata           => open,                           --                      .readdata
			writedata          => open,                           --                      .writedata
			c0                 => open,                           --                    c0.clk
			c1                 => open,                           --                    c1.clk
			c2                 => open,                           --                    c2.clk
			locked             => altpll_0_locked_conduit_export, --        locked_conduit.export
			scandone           => open,                           --           (terminated)
			scandataout        => open,                           --           (terminated)
			c3                 => open,                           --           (terminated)
			c4                 => open,                           --           (terminated)
			areset             => '0',                            --           (terminated)
			phasedone          => open,                           --           (terminated)
			phasecounterselect => "000",                          --           (terminated)
			phaseupdown        => '0',                            --           (terminated)
			phasestep          => '0',                            --           (terminated)
			scanclk            => '0',                            --           (terminated)
			scanclkena         => '0',                            --           (terminated)
			scandata           => '0',                            --           (terminated)
			configupdate       => '0'                             --           (terminated)
		);

	bme280_i2c_0 : component FE_CPLD_BME280_I2C_Reader
		generic map (
			sdo              => '0',
			reads_per_second => 16,
			input_clk        => 50000000
		)
		port map (
			reset_n          => rst_controller_reset_out_reset_ports_inv, --           reset.reset_n
			sys_clk          => clk_clk,                                  --      clock_sink.clk
			bme_output_data  => bme280_i2c_0_bme_output_data,             --      bme_output.data
			bme_output_error => bme280_i2c_0_bme_output_error,            --                .error
			bme_output_valid => bme280_i2c_0_bme_output_valid,            --                .valid
			busy_out         => bme280_i2c_0_control_conduit_busy_out,    -- control_conduit.busy_out
			continuous       => bme280_i2c_0_control_conduit_continuous,  --                .continuous
			enable           => bme280_i2c_0_control_conduit_enable,      --                .enable
			i2c_ack_error    => bme280_i2c_0_i2c_interface_i2c_ack_error, --   I2C_Interface.i2c_ack_error
			i2c_addr         => bme280_i2c_0_i2c_interface_i2c_addr,      --                .i2c_addr
			i2c_busy         => bme280_i2c_0_i2c_interface_i2c_busy,      --                .i2c_busy
			i2c_data_rd      => bme280_i2c_0_i2c_interface_i2c_data_rd,   --                .i2c_data_rd
			i2c_data_wr      => bme280_i2c_0_i2c_interface_i2c_data_wr,   --                .i2c_data_wr
			i2c_ena          => bme280_i2c_0_i2c_interface_i2c_ena,       --                .i2c_ena
			i2c_rw           => bme280_i2c_0_i2c_interface_i2c_rw         --                .i2c_rw
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of cx_system
